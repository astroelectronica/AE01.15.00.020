.title KiCad schematic
V1 /IN 0 AC 1
R1 /IN /H {R}
R3 /H /OUT {R}
C2 /H 0 {CM}
C1 /L /IN {C}
C3 /OUT /L {C}
R2 /L 0 {RM}
.end
